--Lets check if it is saved